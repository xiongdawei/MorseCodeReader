module decoder(
    input      [5:0] morse,
    input      [3:0] sw,
    output reg [3:0] number
);



endmodule