module Counter(
    input            clk,
    input            reset,
    input            enable,
    input            clear,
    output reg [3:0] q
);

// YOU NEED TO EDIT THE ALWAYS BLOCK TO IMPLEMENT THE COUNTER

always @(posedge clk, posedge reset) begin
end

endmodule